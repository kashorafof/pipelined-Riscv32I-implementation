
`ifndef Memory_definitions
`define Memory_definitions

`define Word 2'b00
`define Half 2'b01
`define Byte 2'b10
`define Signed 1'b1
`define Unsigned 1'b0

`define Read 1'b0
`define Write 1'b1
`endif
