`define I_format 3'b000
`define S_format 3'b001
`define B_format 3'b010
`define U_format 3'b011
`define J_format 3'b100
