parameter Word = 2'b00;
parameter Half = 2'b01;
parameter Byte = 2'b10;
parameter Signed = 1'b1;
parameter Unsigned = 1'b0;