module TOP_CPU(
  input wire clk_i, rst_i,
  input wire [31:0] Instr_i,
  
);






endmodule