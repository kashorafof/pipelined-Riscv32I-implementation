parameter I_format = 3'b000;
parameter S_format = 3'b001;
parameter B_format = 3'b010;
parameter U_format = 3'b011;
parameter J_format = 3'b100;
