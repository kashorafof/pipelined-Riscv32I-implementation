parameter ADD = 4'b0000;
parameter SUB = 4'b0001;
parameter SLL = 4'b0010;
parameter SRL = 4'b0011;
parameter SRA = 4'b0100;
parameter XOR = 4'b0101;
parameter AND = 4'b0110;
parameter OR = 4'b0111;
parameter SLT = 4'b1000;
parameter SLTU = 4'b1001;
parameter EQ = 4'b1010;
parameter NE = 4'b1011;
parameter LT = 4'b1100;
parameter GE = 4'b1101;
parameter LTU = 4'b1110;
parameter GEU = 4'b1111;