`ifndef alu_definitions
`define alu_definitions

`define ADD 4'b0000
`define SUB 4'b0001
`define SLL 4'b0010
`define SRL 4'b0011
`define SRA 4'b0100
`define XOR 4'b0101
`define AND 4'b0110
`define OR 4'b0111
`define SLT 4'b1000
`define SLTU 4'b1001

`endif
