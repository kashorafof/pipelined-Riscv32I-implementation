`ifndef Format_definitions
`define Format_definitions

`define I_Format 3'b000
`define S_Format 3'b001
`define B_Format 3'b010
`define U_Format 3'b011
`define J_Format 3'b100
`define R_Format 3'b101

`endif  // Format_definitions
