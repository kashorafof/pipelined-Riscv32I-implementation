`ifndef alu_definitions
`define alu_definitions

`define ADD 4'b0000
`define SUB 4'b0001
`define SLL 4'b0010
`define SRL 4'b0011
`define SRA 4'b0100
`define XOR 4'b0101
`define AND 4'b0110
`define OR 4'b0111
`define SLT 4'b1000
`define SLTU 4'b1001
`define EQ 4'b1010
`define NE 4'b1011
`define LT 4'b1100
`define GE 4'b1101
`define LTU 4'b1110
`define GEU 4'b1111

`endif
